magic
tech sky130A
magscale 1 2
timestamp 1711885615
<< error_s >>
rect 5650 7500 5708 7506
rect 5650 7466 5662 7500
rect 5650 7460 5708 7466
rect 5650 7172 5708 7178
rect 5650 7138 5662 7172
rect 5650 7132 5708 7138
rect 5636 5848 5694 5854
rect 5636 5814 5648 5848
rect 5636 5808 5694 5814
rect 5636 5538 5694 5544
rect 5636 5504 5648 5538
rect 5636 5498 5694 5504
<< metal1 >>
rect 132 14754 388 14998
rect 156 14752 356 14754
rect -1780 8094 -1516 8106
rect -1780 7894 8912 8094
rect -1780 7844 -1516 7894
rect -1744 6762 -1480 6788
rect -1744 6570 8848 6762
rect -1744 6562 -1260 6570
rect -506 6562 -436 6570
rect -1744 6526 -1480 6562
rect 5302 -588 5366 -586
rect 5276 -796 5492 -588
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1711880980
transform 1 0 6664 0 1 11124
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1711880980
transform 1 0 5665 0 1 5676
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1711880980
transform 1 0 5679 0 1 7319
box -211 -319 211 319
use sky130_fd_pr__res_high_po_0p35_TTBX7G  XR1
timestamp 1711880980
transform 1 0 148 0 1 7129
box -201 -6582 201 6582
<< labels >>
flabel metal1 -1780 7844 -1516 8106 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
flabel metal1 -1744 6526 -1480 6788 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 5276 -796 5492 -588 0 FreeSans 1600 0 0 0 out
port 8 nsew
flabel metal1 132 14754 388 14998 0 FreeSans 1600 0 0 0 in
port 6 nsew
<< end >>
