VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_magic_challenge
  CLASS BLOCK ;
  FOREIGN tt_um_magic_challenge ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 154.870 224.760 155.170 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 158.550 224.760 158.850 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.190 224.760 151.490 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 156.560 0.000 157.160 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 134.480 0.000 135.080 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 112.400 0.000 113.000 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 90.320 0.000 90.920 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 68.240 0.000 68.840 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 46.160 0.000 46.760 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 24.080 0.000 24.680 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 2.000 0.000 2.600 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met4 ;
        RECT 147.510 224.760 147.810 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.279000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 140.150 224.760 140.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.470 224.760 136.770 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 129.110 224.760 129.410 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.070 224.760 118.370 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.030 224.760 107.330 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.990 224.760 96.290 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 29.750 224.760 30.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 22.390 224.760 22.690 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 18.710 224.760 19.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 11.350 224.760 11.650 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 7.670 224.760 7.970 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 3.990 224.760 4.290 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 51.830 224.760 52.130 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 40.790 224.760 41.090 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.546900 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.950 224.760 85.250 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 73.910 224.760 74.210 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 62.870 224.760 63.170 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 49.000 5.000 50.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 113.170 208.040 114.010 208.120 ;
        RECT 117.300 208.040 119.120 208.435 ;
        RECT 113.170 206.650 119.120 208.040 ;
        RECT 113.170 206.515 114.010 206.650 ;
        RECT 117.300 206.575 119.120 206.650 ;
      LAYER pwell ;
        RECT 113.375 205.400 113.805 206.185 ;
        RECT 117.510 205.160 118.880 206.155 ;
        RECT 117.490 204.915 118.930 205.160 ;
      LAYER li1 ;
        RECT 117.490 208.160 118.930 208.330 ;
        RECT 113.360 207.845 113.820 208.015 ;
        RECT 113.445 206.680 113.735 207.845 ;
        RECT 117.595 206.735 117.925 208.160 ;
        RECT 117.595 206.405 117.925 206.465 ;
        RECT 116.205 206.215 117.925 206.405 ;
        RECT 113.445 205.295 113.735 206.020 ;
        RECT 116.205 205.955 116.395 206.215 ;
        RECT 117.595 206.095 117.925 206.215 ;
        RECT 118.095 206.095 118.325 207.895 ;
        RECT 118.495 206.735 118.825 208.160 ;
        RECT 118.495 206.460 118.825 206.465 ;
        RECT 118.495 206.160 120.700 206.460 ;
        RECT 118.495 206.095 118.825 206.160 ;
        RECT 118.155 205.925 118.325 206.095 ;
        RECT 113.360 205.125 113.820 205.295 ;
        RECT 117.620 205.000 117.950 205.925 ;
        RECT 118.155 205.755 118.770 205.925 ;
        RECT 118.440 205.265 118.770 205.755 ;
        RECT 117.490 204.830 118.930 205.000 ;
        RECT 116.250 203.950 116.990 204.070 ;
        RECT 113.965 203.255 116.990 203.950 ;
        RECT 116.250 203.150 116.990 203.255 ;
      LAYER mcon ;
        RECT 117.645 208.160 117.815 208.330 ;
        RECT 118.125 208.160 118.295 208.330 ;
        RECT 118.605 208.160 118.775 208.330 ;
        RECT 113.505 207.845 113.675 208.015 ;
        RECT 118.155 207.120 118.325 207.290 ;
        RECT 116.215 205.965 116.385 206.135 ;
        RECT 120.430 206.190 120.670 206.430 ;
        RECT 113.505 205.125 113.675 205.295 ;
        RECT 117.645 204.830 117.815 205.000 ;
        RECT 118.125 204.830 118.295 205.000 ;
        RECT 118.605 204.830 118.775 205.000 ;
        RECT 113.995 203.285 114.630 203.920 ;
      LAYER met1 ;
        RECT 104.570 208.550 106.070 209.050 ;
        RECT 104.570 207.995 119.365 208.550 ;
        RECT 104.570 207.490 106.070 207.995 ;
        RECT 113.360 207.690 113.820 207.995 ;
        RECT 116.420 207.300 117.150 207.350 ;
        RECT 118.095 207.300 118.385 207.320 ;
        RECT 116.420 207.105 118.385 207.300 ;
        RECT 116.420 207.050 117.150 207.105 ;
        RECT 118.095 207.090 118.385 207.105 ;
        RECT 115.620 206.580 115.980 206.880 ;
        RECT 115.650 206.390 115.950 206.580 ;
        RECT 115.725 206.145 115.915 206.390 ;
        RECT 116.185 206.145 116.415 206.195 ;
        RECT 120.370 206.160 120.730 206.460 ;
        RECT 115.725 205.955 116.415 206.145 ;
        RECT 116.185 205.905 116.415 205.955 ;
        RECT 104.000 205.110 105.430 205.540 ;
        RECT 113.360 205.110 113.820 205.450 ;
        RECT 120.400 205.370 120.700 206.160 ;
        RECT 117.490 205.110 118.930 205.160 ;
        RECT 104.000 204.415 119.045 205.110 ;
        RECT 120.370 205.070 120.730 205.370 ;
        RECT 104.000 203.980 105.430 204.415 ;
        RECT 113.965 203.950 114.660 204.415 ;
        RECT 113.935 203.255 114.690 203.950 ;
      LAYER via ;
        RECT 104.570 207.520 106.070 209.020 ;
        RECT 116.450 207.050 116.750 207.350 ;
        RECT 115.650 206.580 115.950 206.880 ;
        RECT 104.000 204.010 105.430 205.510 ;
        RECT 120.400 205.070 120.700 205.370 ;
      LAYER met2 ;
        RECT 102.125 209.020 103.575 209.040 ;
        RECT 102.100 207.520 106.100 209.020 ;
        RECT 116.450 207.830 116.750 207.840 ;
        RECT 115.650 207.630 115.950 207.640 ;
        RECT 102.125 207.500 103.575 207.520 ;
        RECT 115.615 207.350 115.985 207.630 ;
        RECT 116.415 207.550 116.785 207.830 ;
        RECT 115.650 206.550 115.950 207.350 ;
        RECT 116.450 207.020 116.750 207.550 ;
        RECT 103.930 204.565 105.460 205.510 ;
        RECT 120.400 205.370 120.700 205.400 ;
        RECT 121.040 205.370 121.320 205.405 ;
        RECT 120.400 205.070 121.330 205.370 ;
        RECT 120.400 205.040 120.700 205.070 ;
        RECT 121.040 205.035 121.320 205.070 ;
        RECT 103.910 204.010 105.460 204.565 ;
        RECT 103.910 203.115 105.450 204.010 ;
        RECT 103.930 203.090 105.430 203.115 ;
      LAYER via2 ;
        RECT 102.125 207.545 103.575 208.995 ;
        RECT 115.660 207.350 115.940 207.630 ;
        RECT 116.460 207.550 116.740 207.830 ;
        RECT 121.040 205.080 121.320 205.360 ;
        RECT 103.955 203.115 105.405 204.565 ;
      LAYER met3 ;
        RECT 115.610 209.270 115.990 209.590 ;
        RECT 36.885 209.020 38.375 209.045 ;
        RECT 36.880 207.520 103.630 209.020 ;
        RECT 115.650 207.655 115.950 209.270 ;
        RECT 116.410 208.330 116.790 208.650 ;
        RECT 116.450 207.855 116.750 208.330 ;
        RECT 36.885 207.495 38.375 207.520 ;
        RECT 115.635 207.325 115.965 207.655 ;
        RECT 116.435 207.525 116.765 207.855 ;
        RECT 120.990 205.750 121.370 206.070 ;
        RECT 121.030 205.385 121.330 205.750 ;
        RECT 121.015 205.055 121.345 205.385 ;
        RECT 103.930 202.895 105.430 204.590 ;
        RECT 103.905 201.405 105.455 202.895 ;
        RECT 103.930 201.400 105.430 201.405 ;
      LAYER via3 ;
        RECT 115.640 209.270 115.960 209.590 ;
        RECT 36.885 207.525 38.375 209.015 ;
        RECT 116.440 208.330 116.760 208.650 ;
        RECT 121.020 205.750 121.340 206.070 ;
        RECT 103.935 201.405 105.425 202.895 ;
      LAYER met4 ;
        RECT 88.630 214.210 88.930 224.760 ;
        RECT 88.630 213.910 117.050 214.210 ;
        RECT 116.700 211.040 117.000 213.910 ;
        RECT 143.830 212.090 144.130 224.760 ;
        RECT 118.270 211.790 144.130 212.090 ;
        RECT 114.750 210.740 117.000 211.040 ;
        RECT 2.500 207.520 38.380 209.020 ;
        RECT 114.750 208.640 115.050 210.740 ;
        RECT 115.635 209.580 115.965 209.595 ;
        RECT 118.300 209.580 118.600 211.790 ;
        RECT 143.830 211.720 144.130 211.790 ;
        RECT 147.510 209.720 147.810 224.760 ;
        RECT 115.635 209.280 118.600 209.580 ;
        RECT 121.030 209.420 147.810 209.720 ;
        RECT 115.635 209.265 115.965 209.280 ;
        RECT 116.435 208.640 116.765 208.655 ;
        RECT 114.750 208.340 116.765 208.640 ;
        RECT 114.750 208.330 115.050 208.340 ;
        RECT 116.435 208.325 116.765 208.340 ;
        RECT 121.030 206.075 121.330 209.420 ;
        RECT 121.015 205.745 121.345 206.075 ;
        RECT 50.500 201.400 105.430 202.900 ;
  END
END tt_um_magic_challenge
END LIBRARY

