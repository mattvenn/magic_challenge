magic
tech sky130A
magscale 1 2
timestamp 1711885285
<< metal1 >>
rect 24704 18960 24824 18966
rect 24472 18840 24704 18960
rect 24472 17750 24592 18840
rect 24704 18834 24824 18840
rect 19398 11126 19698 11132
rect 19698 10826 22736 11126
rect 19398 10820 19698 10826
rect 19220 9492 19226 9792
rect 19526 9492 22678 9792
rect 28242 2346 28362 2352
rect 28362 2226 29758 2346
rect 28242 2220 28362 2226
<< via1 >>
rect 24704 18840 24824 18960
rect 19398 10826 19698 11126
rect 19226 9492 19526 9792
rect 28242 2226 28362 2346
<< metal2 >>
rect 26113 18960 26223 18964
rect 24698 18840 24704 18960
rect 24824 18955 26228 18960
rect 24824 18845 26113 18955
rect 26223 18845 26228 18955
rect 24824 18840 26228 18845
rect 26113 18836 26223 18840
rect 17443 11126 17733 11130
rect 17438 11121 19398 11126
rect 17438 10831 17443 11121
rect 17733 10831 19398 11121
rect 17438 10826 19398 10831
rect 19698 10826 19704 11126
rect 17443 10822 17733 10826
rect 17415 9792 17705 9796
rect 19226 9792 19526 9798
rect 17410 9787 19226 9792
rect 17410 9497 17415 9787
rect 17705 9497 19226 9787
rect 17410 9492 19226 9497
rect 17415 9488 17705 9492
rect 19226 9486 19526 9492
rect 27469 2346 27579 2350
rect 27464 2341 28242 2346
rect 27464 2231 27469 2341
rect 27579 2231 28242 2341
rect 27464 2226 28242 2231
rect 28362 2226 28368 2346
rect 27469 2222 27579 2226
<< via2 >>
rect 26113 18845 26223 18955
rect 17443 10831 17733 11121
rect 17415 9497 17705 9787
rect 27469 2231 27579 2341
<< metal3 >>
rect 28487 18960 28605 18965
rect 26108 18959 28606 18960
rect 26108 18955 28487 18959
rect 26108 18845 26113 18955
rect 26223 18845 28487 18955
rect 26108 18841 28487 18845
rect 28605 18841 28606 18959
rect 26108 18840 28606 18841
rect 28487 18835 28605 18840
rect 5229 11126 5527 11131
rect 5228 11125 17738 11126
rect 5228 10827 5229 11125
rect 5527 11121 17738 11125
rect 5527 10831 17443 11121
rect 17733 10831 17738 11121
rect 5527 10827 17738 10831
rect 5228 10826 17738 10827
rect 5229 10821 5527 10826
rect 14910 9791 17710 9792
rect 14905 9493 14911 9791
rect 15209 9787 17710 9791
rect 15209 9497 17415 9787
rect 17705 9497 17710 9787
rect 15209 9493 17710 9497
rect 14910 9492 17710 9493
rect 26896 2345 27584 2346
rect 26891 2227 26897 2345
rect 27015 2341 27584 2345
rect 27015 2231 27469 2341
rect 27579 2231 27584 2341
rect 27015 2227 27584 2231
rect 26896 2226 27584 2227
<< via3 >>
rect 28487 18841 28605 18959
rect 5229 10827 5527 11125
rect 14911 9493 15209 9791
rect 26897 2227 27015 2345
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 17726 44952 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 200 11126 500 44152
rect 200 11125 5528 11126
rect 200 10827 5229 11125
rect 5527 10827 5528 11125
rect 200 10826 5528 10827
rect 200 1000 500 10826
rect 9800 9792 10100 44152
rect 28486 18959 37392 18960
rect 28486 18841 28487 18959
rect 28605 18841 37392 18959
rect 28486 18840 37392 18841
rect 9800 9791 15210 9792
rect 9800 9493 14911 9791
rect 15209 9493 15210 9791
rect 9800 9492 15210 9493
rect 9800 1000 10100 9492
rect 26896 2345 27016 2346
rect 26896 2227 26897 2345
rect 27015 2227 27016 2345
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 2227
rect 37272 1366 37392 18840
rect 31312 1246 37392 1366
rect 31312 0 31432 1246
use challenge  challenge_0 ~/work/asic-workshop/shuttle-2404/magic-challenge/mag
timestamp 1711885285
transform 1 0 24307 0 1 2986
box -1780 -796 10180 14998
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
