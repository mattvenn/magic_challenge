magic
tech sky130A
magscale 1 2
timestamp 1710074111
<< pwell >>
rect -199 -1596 199 1596
<< psubdiff >>
rect -163 1526 -67 1560
rect 67 1526 163 1560
rect -163 1464 -129 1526
rect 129 1464 163 1526
rect -163 -1526 -129 -1464
rect 129 -1526 163 -1464
rect -163 -1560 -67 -1526
rect 67 -1560 163 -1526
<< psubdiffcont >>
rect -67 1526 67 1560
rect -163 -1464 -129 1464
rect 129 -1464 163 1464
rect -67 -1560 67 -1526
<< poly >>
rect -33 1414 33 1430
rect -33 1380 -17 1414
rect 17 1380 33 1414
rect -33 1000 33 1380
rect -33 -1380 33 -1000
rect -33 -1414 -17 -1380
rect 17 -1414 33 -1380
rect -33 -1430 33 -1414
<< polycont >>
rect -17 1380 17 1414
rect -17 -1414 17 -1380
<< npolyres >>
rect -33 -1000 33 1000
<< locali >>
rect -163 1526 -67 1560
rect 67 1526 163 1560
rect -163 1464 -129 1526
rect 129 1464 163 1526
rect -33 1380 -17 1414
rect 17 1380 33 1414
rect -33 -1414 -17 -1380
rect 17 -1414 33 -1380
rect -163 -1526 -129 -1464
rect 129 -1526 163 -1464
rect -163 -1560 -67 -1526
rect 67 -1560 163 -1526
<< viali >>
rect -17 1380 17 1414
rect -17 1017 17 1380
rect -17 -1380 17 -1017
rect -17 -1414 17 -1380
<< metal1 >>
rect -23 1414 23 1426
rect -23 1017 -17 1414
rect 17 1017 23 1414
rect -23 1005 23 1017
rect -23 -1017 23 -1005
rect -23 -1414 -17 -1017
rect 17 -1414 23 -1017
rect -23 -1426 23 -1414
<< properties >>
string FIXED_BBOX -146 -1543 146 1543
string gencell sky130_fd_pr__res_generic_po
string library sky130
string parameters w 0.330 l 10 m 1 nx 1 wmin 0.330 lmin 1.650 rho 48.2 val 1.46k dummy 0 dw 0.0 term 0.0 sterm 0.0 caplen 0.4 snake 0 guard 1 glc 1 grc 1 gtc 1 gbc 1 roverlap 0 endcov 100 full_metal 1 hv_guard 0 n_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
