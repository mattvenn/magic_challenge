magic
tech sky130A
magscale 1 2
timestamp 1727432336
<< viali >>
rect 5640 7564 5732 7606
rect 264 6598 322 6744
rect 5600 5914 5732 5952
<< metal1 >>
rect 132 14754 388 14998
rect 156 14752 356 14754
rect -1780 8094 -1516 8106
rect -1780 7894 8912 8094
rect -1780 7844 -1516 7894
rect 5322 7384 5448 7894
rect 5628 7642 5742 7894
rect 5620 7606 5750 7642
rect 5620 7564 5640 7606
rect 5732 7564 5750 7606
rect 5620 7550 5750 7564
rect 5642 7458 6614 7510
rect 5322 7258 5652 7384
rect 5698 7270 6074 7386
rect 6190 7270 6196 7386
rect 6562 7324 6614 7458
rect 7222 7324 7386 7330
rect 6562 7182 7222 7324
rect 5650 7160 7222 7182
rect 5650 7130 6614 7160
rect 7222 7154 7386 7160
rect 6558 6988 6610 7130
rect 6558 6930 6610 6936
rect -1744 6762 -1480 6788
rect -1744 6744 8848 6762
rect -1744 6598 264 6744
rect 322 6598 8848 6744
rect -1744 6570 8848 6598
rect -1744 6562 -1260 6570
rect -506 6562 -436 6570
rect -1744 6526 -1480 6562
rect 5326 5734 5434 6570
rect 5582 5952 5754 6570
rect 5582 5914 5600 5952
rect 5732 5914 5754 5952
rect 5582 5900 5754 5914
rect 6558 6366 6610 6372
rect 5626 5808 6280 5860
rect 5326 5626 5644 5734
rect 5688 5618 6074 5734
rect 6190 5618 6196 5734
rect 6224 5708 6276 5808
rect 6558 5708 6610 6314
rect 6224 5656 6610 5708
rect 6224 5546 6276 5656
rect 5626 5494 6276 5546
rect 6296 4890 6302 5098
rect 6510 4890 6516 5098
rect 6302 3046 6510 4890
rect 5276 2838 6510 3046
rect 1034 2510 1194 2516
rect 1034 994 1194 2350
rect 72 834 1194 994
rect 5276 -588 5484 2838
rect 5276 -796 5492 -588
<< via1 >>
rect 6074 7270 6190 7386
rect 7222 7160 7386 7324
rect 6558 6936 6610 6988
rect 6558 6314 6610 6366
rect 6074 5618 6190 5734
rect 6302 4890 6510 5098
rect 1034 2350 1194 2510
<< metal2 >>
rect 1034 10426 1556 10586
rect 1716 10426 1725 10586
rect 1034 2510 1194 10426
rect 7222 7559 7386 7564
rect 7218 7405 7227 7559
rect 7381 7405 7390 7559
rect 6074 7386 6190 7392
rect 7222 7324 7386 7405
rect 6074 6180 6190 7270
rect 7216 7160 7222 7324
rect 7386 7160 7392 7324
rect 6552 6936 6558 6988
rect 6610 6936 6616 6988
rect 6558 6366 6610 6936
rect 6552 6314 6558 6366
rect 6610 6314 6616 6366
rect 6074 5972 6510 6180
rect 6074 5734 6190 5972
rect 6074 5612 6190 5618
rect 6302 5098 6510 5972
rect 6302 4884 6510 4890
rect 1028 2350 1034 2510
rect 1194 2350 1200 2510
<< via2 >>
rect 1556 10426 1716 10586
rect 7227 7405 7381 7559
<< metal3 >>
rect 1551 10586 1721 10591
rect 1551 10426 1556 10586
rect 1716 10426 2324 10586
rect 2484 10426 2490 10586
rect 1551 10421 1721 10426
rect 7222 7789 7386 7790
rect 7217 7627 7223 7789
rect 7385 7627 7391 7789
rect 7222 7559 7386 7627
rect 7222 7405 7227 7559
rect 7381 7405 7386 7559
rect 7222 7400 7386 7405
<< via3 >>
rect 2324 10426 2484 10586
rect 7223 7627 7385 7789
<< metal4 >>
rect 2323 10586 2485 10587
rect 2323 10426 2324 10586
rect 2484 10426 5404 10586
rect 2323 10425 2485 10426
rect 8734 8910 8898 9790
rect 7222 8746 8898 8910
rect 7222 7789 7386 8746
rect 7222 7627 7223 7789
rect 7385 7627 7386 7789
rect 7222 7626 7386 7627
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1711880980
transform 1 0 6664 0 1 11124
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1727432252
transform 1 0 5665 0 1 5676
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1727432252
transform 1 0 5679 0 1 7319
box -211 -319 211 319
use sky130_fd_pr__res_high_po_0p35_TTBX7G  XR1
timestamp 1711880980
transform 1 0 148 0 1 7129
box -201 -6582 201 6582
<< labels >>
flabel metal1 -1780 7844 -1516 8106 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
flabel metal1 -1744 6526 -1480 6788 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 5276 -796 5492 -588 0 FreeSans 1600 0 0 0 out
port 8 nsew
flabel metal1 132 14754 388 14998 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel metal2 1034 2510 1194 10586 0 FreeSans 1600 0 0 0 tocap
flabel metal4 7222 7789 7386 8910 0 FreeSans 1600 0 0 0 gate
<< end >>
