magic
tech sky130A
magscale 1 2
timestamp 1710086986
<< nwell >>
rect 22652 41330 23802 41608
<< psubdiff >>
rect 23250 40798 23398 40822
rect 23250 40622 23398 40646
<< psubdiffcont >>
rect 23250 40646 23398 40798
<< locali >>
rect 23706 41286 24140 41292
rect 23241 41243 23573 41281
rect 23241 41227 23279 41243
rect 23706 41238 24086 41286
rect 24134 41238 24140 41286
rect 23706 41232 24140 41238
rect 23241 41193 23243 41227
rect 23277 41193 23279 41227
rect 23241 41191 23279 41193
rect 23250 40798 23398 40814
rect 22793 40784 23250 40790
rect 22793 40657 22799 40784
rect 22926 40657 23250 40784
rect 22793 40651 23250 40657
rect 23250 40630 23398 40646
<< viali >>
rect 23631 41424 23665 41458
rect 24086 41238 24134 41286
rect 23243 41193 23277 41227
rect 22799 40657 22926 40784
<< metal1 >>
rect 20914 41804 21214 41810
rect 21214 41599 23873 41710
rect 20914 41498 21214 41504
rect 23284 41410 23290 41470
rect 23350 41460 23430 41470
rect 23619 41460 23677 41464
rect 23350 41458 23677 41460
rect 23350 41424 23631 41458
rect 23665 41424 23677 41458
rect 23350 41421 23677 41424
rect 23350 41410 23430 41421
rect 23619 41418 23677 41421
rect 23124 41316 23130 41376
rect 23190 41316 23196 41376
rect 23130 41278 23190 41316
rect 24074 41286 24146 41292
rect 23145 41229 23183 41278
rect 23237 41229 23283 41239
rect 24074 41238 24086 41286
rect 24134 41238 24146 41286
rect 24074 41232 24146 41238
rect 23145 41227 23283 41229
rect 23145 41193 23243 41227
rect 23277 41193 23283 41227
rect 23145 41191 23283 41193
rect 23237 41181 23283 41191
rect 20800 41102 21086 41108
rect 24080 41074 24140 41232
rect 21086 40883 23809 41022
rect 24074 41014 24080 41074
rect 24140 41014 24146 41074
rect 20800 40796 21086 40802
rect 22793 40790 22932 40883
rect 22787 40784 22938 40790
rect 22787 40657 22799 40784
rect 22926 40657 22938 40784
rect 22787 40651 22938 40657
rect 27790 4476 27916 4484
rect 27786 4356 28862 4476
rect 28742 4316 28862 4356
rect 29784 4316 29904 4322
rect 28742 4196 29784 4316
rect 29784 4190 29904 4196
rect 26896 1730 27926 1850
rect 26896 1620 27016 1730
rect 26890 1500 26896 1620
rect 27016 1500 27022 1620
<< via1 >>
rect 20914 41504 21214 41804
rect 23290 41410 23350 41470
rect 23130 41316 23190 41376
rect 20800 40802 21086 41102
rect 24080 41014 24140 41074
rect 29784 4196 29904 4316
rect 26896 1500 27016 1620
<< metal2 >>
rect 20425 41804 20715 41808
rect 20420 41799 20914 41804
rect 20420 41509 20425 41799
rect 20715 41509 20914 41799
rect 20420 41504 20914 41509
rect 21214 41504 21220 41804
rect 23290 41566 23350 41568
rect 23130 41526 23190 41528
rect 20425 41500 20715 41504
rect 23123 41470 23132 41526
rect 23188 41470 23197 41526
rect 23283 41510 23292 41566
rect 23348 41510 23357 41566
rect 23290 41470 23350 41510
rect 23130 41376 23190 41470
rect 23290 41404 23350 41410
rect 23130 41310 23190 41316
rect 20786 40913 20800 41102
rect 20782 40623 20791 40913
rect 21086 40802 21092 41102
rect 24080 41074 24140 41080
rect 24208 41074 24264 41081
rect 24140 41072 24266 41074
rect 24140 41016 24208 41072
rect 24264 41016 24266 41072
rect 24140 41014 24266 41016
rect 24080 41008 24140 41014
rect 24208 41007 24264 41014
rect 21081 40623 21090 40802
rect 20786 40618 21086 40623
rect 30293 4316 30403 4320
rect 29778 4196 29784 4316
rect 29904 4311 30408 4316
rect 29904 4201 30293 4311
rect 30403 4201 30408 4311
rect 29904 4196 30408 4201
rect 30293 4192 30403 4196
rect 26896 1620 27016 1626
rect 26896 1055 27016 1500
rect 26892 945 26901 1055
rect 27011 945 27020 1055
rect 26896 940 27016 945
<< via2 >>
rect 20425 41509 20715 41799
rect 23132 41470 23188 41526
rect 23292 41510 23348 41566
rect 20791 40802 20800 40913
rect 20800 40802 21081 40913
rect 24208 41016 24264 41072
rect 20791 40623 21081 40802
rect 30293 4201 30403 4311
rect 26901 945 27011 1055
<< metal3 >>
rect 23122 41854 23128 41918
rect 23192 41854 23198 41918
rect 7377 41804 7675 41809
rect 7376 41803 20726 41804
rect 7376 41505 7377 41803
rect 7675 41799 20726 41803
rect 7675 41509 20425 41799
rect 20715 41509 20726 41799
rect 23130 41531 23190 41854
rect 23282 41666 23288 41730
rect 23352 41666 23358 41730
rect 23290 41571 23350 41666
rect 23287 41566 23353 41571
rect 7675 41505 20726 41509
rect 7376 41504 20726 41505
rect 23127 41526 23193 41531
rect 7377 41499 7675 41504
rect 23127 41470 23132 41526
rect 23188 41470 23193 41526
rect 23287 41510 23292 41566
rect 23348 41510 23353 41566
rect 23287 41505 23353 41510
rect 23127 41465 23193 41470
rect 24198 41150 24204 41214
rect 24268 41150 24274 41214
rect 24206 41077 24266 41150
rect 24203 41072 24269 41077
rect 24203 41016 24208 41072
rect 24264 41016 24269 41072
rect 24203 41011 24269 41016
rect 20786 40913 21086 40918
rect 20786 40623 20791 40913
rect 21081 40623 21086 40913
rect 20786 40579 21086 40623
rect 20781 40281 20787 40579
rect 21085 40281 21091 40579
rect 20786 40280 21086 40281
rect 31313 4316 31431 4321
rect 30288 4315 31432 4316
rect 30288 4311 31313 4315
rect 30288 4201 30293 4311
rect 30403 4201 31313 4311
rect 30288 4197 31313 4201
rect 31431 4197 31432 4315
rect 30288 4196 31432 4197
rect 31313 4191 31431 4196
rect 26896 1055 27016 1060
rect 26896 945 26901 1055
rect 27011 945 27016 1055
rect 26896 839 27016 945
rect 26891 721 26897 839
rect 27015 721 27021 839
rect 26896 720 27016 721
<< via3 >>
rect 23128 41854 23192 41918
rect 7377 41505 7675 41803
rect 23288 41666 23352 41730
rect 24204 41150 24268 41214
rect 20787 40281 21085 40579
rect 31313 4197 31431 4315
rect 26897 721 27015 839
<< metal4 >>
rect 798 44952 858 45152
rect 1534 44952 1594 45152
rect 2270 44952 2330 45152
rect 3006 44952 3066 45152
rect 3742 44952 3802 45152
rect 4478 44952 4538 45152
rect 5214 44952 5274 45152
rect 5950 44952 6010 45152
rect 6686 44952 6746 45152
rect 7422 44952 7482 45152
rect 8158 44952 8218 45152
rect 8894 44952 8954 45152
rect 9630 44952 9690 45152
rect 10366 44952 10426 45152
rect 11102 44952 11162 45152
rect 11838 44952 11898 45152
rect 12574 44952 12634 45152
rect 13310 44952 13370 45152
rect 14046 44952 14106 45152
rect 14782 44952 14842 45152
rect 15518 44952 15578 45152
rect 16254 44952 16314 45152
rect 16990 44952 17050 45152
rect 200 41804 500 44152
rect 200 41803 7676 41804
rect 200 41505 7377 41803
rect 7675 41505 7676 41803
rect 200 41504 7676 41505
rect 200 1000 500 41504
rect 9800 40580 10100 44152
rect 17726 42842 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 17726 42782 23410 42842
rect 23340 42208 23400 42782
rect 28766 42418 28826 45152
rect 23654 42358 28826 42418
rect 22950 42148 23400 42208
rect 22950 41728 23010 42148
rect 23127 41918 23193 41919
rect 23127 41854 23128 41918
rect 23192 41916 23193 41918
rect 23660 41916 23720 42358
rect 28766 42344 28826 42358
rect 29502 41944 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 23192 41856 23720 41916
rect 24206 41884 29562 41944
rect 23192 41854 23193 41856
rect 23127 41853 23193 41854
rect 23287 41730 23353 41731
rect 23287 41728 23288 41730
rect 22950 41668 23288 41728
rect 22950 41666 23010 41668
rect 23287 41666 23288 41668
rect 23352 41666 23353 41730
rect 23287 41665 23353 41666
rect 24206 41215 24266 41884
rect 24203 41214 24269 41215
rect 24203 41150 24204 41214
rect 24268 41150 24269 41214
rect 24203 41149 24269 41150
rect 9800 40579 21086 40580
rect 9800 40281 20787 40579
rect 21085 40281 21086 40579
rect 9800 40280 21086 40281
rect 9800 1000 10100 40280
rect 31312 4315 31432 4316
rect 31312 4197 31313 4315
rect 31431 4197 31432 4315
rect 26896 839 27016 840
rect 26896 721 26897 839
rect 27015 721 27016 839
rect 400 0 520 200
rect 4816 0 4936 200
rect 9232 0 9352 200
rect 13648 0 13768 200
rect 18064 0 18184 200
rect 22480 0 22600 200
rect 26896 0 27016 721
rect 31312 0 31432 4197
use sky130_fd_io__nand2_1  sky130_fd_io__nand2_1_0 $PDKPATH/libs.ref/sky130_fd_io/mag
timestamp 1676037725
transform 1 0 23498 0 1 40983
box -38 -49 326 715
use cells/sky130_fd_pr__res_high_po_0p35_SKZWQ5  sky130_fd_pr__res_high_po_0p35_SKZWQ5_0
timestamp 1710086986
transform 1 0 27797 0 1 2984
box -201 -1598 201 1598
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1685868990
transform 1 0 22672 0 1 41042
box -38 -48 130 592
<< labels >>
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31312 0 31432 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26896 0 27016 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22480 0 22600 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18064 0 18184 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 13648 0 13768 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 9232 0 9352 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4816 0 4936 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 400 0 520 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VPWR
port 51 nsew power bidirectional
flabel metal4 9800 1000 10100 44152 1 FreeSans 2 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
