magic
tech sky130A
magscale 1 2
timestamp 1711885285
<< viali >>
rect 5636 7562 5722 7608
rect 258 6594 326 6740
rect 5632 5916 5696 5952
<< metal1 >>
rect 132 14754 388 14998
rect 156 14730 356 14754
rect 173 14207 339 14730
rect -499 14041 339 14207
rect -498 13370 -334 14041
rect -498 13206 236 13370
rect -1780 8094 -1516 8106
rect -1780 7894 10132 8094
rect -1780 7844 -1516 7894
rect 5280 7362 5364 7894
rect 5610 7608 5756 7894
rect 5610 7562 5636 7608
rect 5722 7562 5756 7608
rect 5610 7552 5756 7562
rect 5638 7452 6004 7504
rect 6056 7452 6062 7504
rect 5280 7298 5650 7362
rect 6764 7352 6828 7358
rect 5284 7290 5650 7298
rect 5710 7288 6764 7352
rect 6764 7282 6828 7288
rect 5924 7174 6004 7176
rect 5648 7124 6004 7174
rect 6056 7124 6062 7176
rect 5648 7122 5970 7124
rect -1744 6762 -1480 6788
rect -1744 6740 10180 6762
rect -1744 6594 258 6740
rect 326 6594 10180 6740
rect -1744 6570 10180 6594
rect -1744 6562 -1260 6570
rect -506 6562 10180 6570
rect -1744 6526 -1480 6562
rect 5282 5714 5386 6562
rect 5594 5952 5752 6562
rect 5594 5916 5632 5952
rect 5696 5916 5752 5952
rect 5594 5910 5752 5916
rect 5638 5846 5696 5848
rect 6092 5846 6098 5855
rect 5638 5812 6098 5846
rect 5638 5808 5696 5812
rect 6092 5803 6098 5812
rect 6150 5803 6156 5855
rect 5282 5664 5636 5714
rect 5696 5710 6012 5726
rect 5696 5668 6764 5710
rect 5320 5656 5636 5664
rect 5932 5646 6764 5668
rect 6828 5646 6834 5710
rect 1258 5263 1264 5573
rect 1574 5263 1580 5573
rect 6098 5544 6150 5550
rect 5963 5533 6098 5535
rect 5651 5501 6098 5533
rect 5651 5499 6042 5501
rect 6098 5486 6150 5492
rect 1264 1084 1574 5263
rect 90 774 1574 1084
rect 5296 102 5302 166
rect 5366 102 5372 166
rect 5302 -588 5366 102
rect 5276 -796 5492 -588
<< via1 >>
rect 6004 7452 6056 7504
rect 6764 7288 6828 7352
rect 6004 7124 6056 7176
rect 6098 5803 6150 5855
rect 6764 5646 6828 5710
rect 1264 5263 1574 5573
rect 6098 5492 6150 5544
rect 5302 102 5366 166
<< metal2 >>
rect 2337 12941 2647 13067
rect 2328 12631 2337 12941
rect 2647 12631 2656 12941
rect 2337 11387 2647 12631
rect 1264 11077 2672 11387
rect 1264 5573 1574 11077
rect 6204 7587 6304 7592
rect 6004 7504 6056 7510
rect 6200 7498 6209 7587
rect 6056 7497 6209 7498
rect 6299 7497 6308 7587
rect 6056 7452 6304 7497
rect 6004 7442 6304 7452
rect 6004 7281 6056 7442
rect 6204 7420 6304 7442
rect 6758 7288 6764 7352
rect 6828 7288 6834 7352
rect 6004 7247 6445 7281
rect 6004 7176 6056 7247
rect 6004 7118 6056 7124
rect 6098 5855 6150 5861
rect 6098 5797 6150 5803
rect 6107 5709 6141 5797
rect 6411 5709 6445 7247
rect 6107 5675 6445 5709
rect 6764 6052 6828 7288
rect 6764 5988 7064 6052
rect 6764 5710 6828 5988
rect 6107 5544 6141 5675
rect 6764 5640 6828 5646
rect 6092 5492 6098 5544
rect 6150 5492 6156 5544
rect 1264 5257 1574 5263
rect 7000 686 7064 5988
rect 5302 622 7064 686
rect 5302 166 5366 622
rect 5302 96 5366 102
<< via2 >>
rect 2337 12631 2647 12941
rect 6209 7497 6299 7587
<< metal3 >>
rect 3342 13509 3348 13819
rect 3658 13509 3664 13819
rect 2332 12941 2652 12946
rect 3348 12941 3658 13509
rect 2332 12631 2337 12941
rect 2647 12631 3658 12941
rect 2332 12626 2652 12631
rect 6204 7727 6304 7728
rect 6199 7629 6205 7727
rect 6303 7629 6309 7727
rect 6204 7587 6304 7629
rect 6204 7497 6209 7587
rect 6299 7497 6304 7587
rect 6204 7492 6304 7497
<< via3 >>
rect 3348 13509 3658 13819
rect 6205 7629 6303 7727
<< metal4 >>
rect 3347 13819 3659 13820
rect 5654 13819 6768 13944
rect 3347 13509 3348 13819
rect 3658 13509 6768 13819
rect 3347 13508 3659 13509
rect 5654 11422 6768 13509
rect 8696 12781 9030 12830
rect 8696 12547 9387 12781
rect 8696 12098 9030 12547
rect 9153 8710 9387 12547
rect 8746 8546 9387 8710
rect 6166 8476 9387 8546
rect 6166 8370 8980 8476
rect 6204 7727 6304 8370
rect 8746 8341 8980 8370
rect 6204 7629 6205 7727
rect 6303 7629 6304 7727
rect 6204 7628 6304 7629
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1711880980
transform 1 0 6664 0 1 11124
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1711880980
transform 1 0 5665 0 1 5676
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1711880980
transform 1 0 5679 0 1 7319
box -211 -319 211 319
use sky130_fd_pr__res_high_po_0p35_TTBX7G  XR1
timestamp 1711880980
transform 1 0 148 0 1 7129
box -201 -6582 201 6582
<< labels >>
flabel metal1 1264 774 1574 5263 0 FreeSans 1600 0 0 0 tocap
flabel metal4 6166 8370 8980 8546 0 FreeSans 1600 0 0 0 gate
flabel metal1 -1780 7844 -1516 8106 0 FreeSans 1600 0 0 0 vdd
port 4 nsew
flabel metal1 -1744 6526 -1480 6788 0 FreeSans 1600 0 0 0 vss
port 5 nsew
flabel metal1 5276 -796 5492 -588 0 FreeSans 1600 0 0 0 out
port 8 nsew
flabel metal1 132 14754 388 14998 0 FreeSans 1600 0 0 0 in
port 6 nsew
<< end >>
